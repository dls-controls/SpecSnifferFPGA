library ieee;
use ieee.std_logic_1164.all;
package spec_defines is
constant FPGA_VERSION: std_logic_vector(15 downto 0)   := X"10_02";
end spec_defines;
