library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity generic_sprom is
    port (
        clk_i : in std_logic;
        addr_i : in unsigned(9 downto 0);
        dat_o : out std_logic_vector(31 downto 0)
    );
end;

architecture rtl of generic_sprom is
    type lookup_t is array(0 to 1023) of std_logic_vector(31 downto 0);
    signal table : lookup_t := (
        X"00000000",
        X"00000001",
        X"00000002",
        X"00000003",
        X"00000004",
        X"00000005",
        X"00000006",
        X"00000007",
        X"00000008",
        X"00000009",
        X"0000000a",
        X"0000000b",
        X"0000000c",
        X"0000000d",
        X"0000000e",
        X"0000000f",
        X"00000010",
        X"00000011",
        X"00000012",
        X"00000013",
        X"00000014",
        X"00000015",
        X"00000016",
        X"00000017",
        X"00000018",
        X"00000019",
        X"0000001a",
        X"0000001b",
        X"0000001c",
        X"0000001d",
        X"0000001e",
        X"0000001f",
        X"00000020",
        X"00000021",
        X"00000022",
        X"00000023",
        X"00000024",
        X"00000025",
        X"00000026",
        X"00000027",
        X"00000028",
        X"00000029",
        X"0000002a",
        X"0000002b",
        X"0000002c",
        X"0000002d",
        X"0000002e",
        X"0000002f",
        X"00000030",
        X"00000031",
        X"00000032",
        X"00000033",
        X"00000034",
        X"00000035",
        X"00000036",
        X"00000037",
        X"00000038",
        X"00000039",
        X"0000003a",
        X"0000003b",
        X"0000003c",
        X"0000003d",
        X"0000003e",
        X"0000003f",
        X"00000040",
        X"00000041",
        X"00000042",
        X"00000043",
        X"00000044",
        X"00000045",
        X"00000046",
        X"00000047",
        X"00000048",
        X"00000049",
        X"0000004a",
        X"0000004b",
        X"0000004c",
        X"0000004d",
        X"0000004e",
        X"0000004f",
        X"00000050",
        X"00000051",
        X"00000052",
        X"00000053",
        X"00000054",
        X"00000055",
        X"00000056",
        X"00000057",
        X"00000058",
        X"00000059",
        X"0000005a",
        X"0000005b",
        X"0000005c",
        X"0000005d",
        X"0000005e",
        X"0000005f",
        X"00000060",
        X"00000061",
        X"00000062",
        X"00000063",
        X"00000064",
        X"00000065",
        X"00000066",
        X"00000067",
        X"00000068",
        X"00000069",
        X"0000006a",
        X"0000006b",
        X"0000006c",
        X"0000006d",
        X"0000006e",
        X"0000006f",
        X"00000070",
        X"00000071",
        X"00000072",
        X"00000073",
        X"00000074",
        X"00000075",
        X"00000076",
        X"00000077",
        X"00000078",
        X"00000079",
        X"0000007a",
        X"0000007b",
        X"0000007c",
        X"0000007d",
        X"0000007e",
        X"0000007f",
        X"00000080",
        X"00000081",
        X"00000082",
        X"00000083",
        X"00000084",
        X"00000085",
        X"00000086",
        X"00000087",
        X"00000088",
        X"00000089",
        X"0000008a",
        X"0000008b",
        X"0000008c",
        X"0000008d",
        X"0000008e",
        X"0000008f",
        X"00000090",
        X"00000091",
        X"00000092",
        X"00000093",
        X"00000094",
        X"00000095",
        X"00000096",
        X"00000097",
        X"00000098",
        X"00000099",
        X"0000009a",
        X"0000009b",
        X"0000009c",
        X"0000009d",
        X"0000009e",
        X"0000009f",
        X"000000a0",
        X"000000a1",
        X"000000a2",
        X"000000a3",
        X"000000a4",
        X"000000a5",
        X"000000a6",
        X"000000a7",
        X"000000a8",
        X"000000a9",
        X"000000aa",
        X"000000ab",
        X"000000ac",
        X"000000ad",
        X"000000ae",
        X"000000af",
        X"000000b0",
        X"000000b1",
        X"000000b2",
        X"000000b3",
        X"000000b4",
        X"000000b5",
        X"000000b6",
        X"000000b7",
        X"000000b8",
        X"000000b9",
        X"000000ba",
        X"000000bb",
        X"000000bc",
        X"000000bd",
        X"000000be",
        X"000000bf",
        X"000000c0",
        X"000000c1",
        X"000000c2",
        X"000000c3",
        X"000000c4",
        X"000000c5",
        X"000000c6",
        X"000000c7",
        X"000000c8",
        X"000000c9",
        X"000000ca",
        X"000000cb",
        X"000000cc",
        X"000000cd",
        X"000000ce",
        X"000000cf",
        X"000000d0",
        X"000000d1",
        X"000000d2",
        X"000000d3",
        X"000000d4",
        X"000000d5",
        X"000000d6",
        X"000000d7",
        X"000000d8",
        X"000000d9",
        X"000000da",
        X"000000db",
        X"000000dc",
        X"000000dd",
        X"000000de",
        X"000000df",
        X"000000e0",
        X"000000e1",
        X"000000e2",
        X"000000e3",
        X"000000e4",
        X"000000e5",
        X"000000e6",
        X"000000e7",
        X"000000e8",
        X"000000e9",
        X"000000ea",
        X"000000eb",
        X"000000ec",
        X"000000ed",
        X"000000ee",
        X"000000ef",
        X"000000f0",
        X"000000f1",
        X"000000f2",
        X"000000f3",
        X"000000f4",
        X"000000f5",
        X"000000f6",
        X"000000f7",
        X"000000f8",
        X"000000f9",
        X"000000fa",
        X"000000fb",
        X"000000fc",
        X"000000fd",
        X"000000fe",
        X"000000ff",
        X"00000100",
        X"00000101",
        X"00000102",
        X"00000103",
        X"00000104",
        X"00000105",
        X"00000106",
        X"00000107",
        X"00000108",
        X"00000109",
        X"0000010a",
        X"0000010b",
        X"0000010c",
        X"0000010d",
        X"0000010e",
        X"0000010f",
        X"00000110",
        X"00000111",
        X"00000112",
        X"00000113",
        X"00000114",
        X"00000115",
        X"00000116",
        X"00000117",
        X"00000118",
        X"00000119",
        X"0000011a",
        X"0000011b",
        X"0000011c",
        X"0000011d",
        X"0000011e",
        X"0000011f",
        X"00000120",
        X"00000121",
        X"00000122",
        X"00000123",
        X"00000124",
        X"00000125",
        X"00000126",
        X"00000127",
        X"00000128",
        X"00000129",
        X"0000012a",
        X"0000012b",
        X"0000012c",
        X"0000012d",
        X"0000012e",
        X"0000012f",
        X"00000130",
        X"00000131",
        X"00000132",
        X"00000133",
        X"00000134",
        X"00000135",
        X"00000136",
        X"00000137",
        X"00000138",
        X"00000139",
        X"0000013a",
        X"0000013b",
        X"0000013c",
        X"0000013d",
        X"0000013e",
        X"0000013f",
        X"00000140",
        X"00000141",
        X"00000142",
        X"00000143",
        X"00000144",
        X"00000145",
        X"00000146",
        X"00000147",
        X"00000148",
        X"00000149",
        X"0000014a",
        X"0000014b",
        X"0000014c",
        X"0000014d",
        X"0000014e",
        X"0000014f",
        X"00000150",
        X"00000151",
        X"00000152",
        X"00000153",
        X"00000154",
        X"00000155",
        X"00000156",
        X"00000157",
        X"00000158",
        X"00000159",
        X"0000015a",
        X"0000015b",
        X"0000015c",
        X"0000015d",
        X"0000015e",
        X"0000015f",
        X"00000160",
        X"00000161",
        X"00000162",
        X"00000163",
        X"00000164",
        X"00000165",
        X"00000166",
        X"00000167",
        X"00000168",
        X"00000169",
        X"0000016a",
        X"0000016b",
        X"0000016c",
        X"0000016d",
        X"0000016e",
        X"0000016f",
        X"00000170",
        X"00000171",
        X"00000172",
        X"00000173",
        X"00000174",
        X"00000175",
        X"00000176",
        X"00000177",
        X"00000178",
        X"00000179",
        X"0000017a",
        X"0000017b",
        X"0000017c",
        X"0000017d",
        X"0000017e",
        X"0000017f",
        X"00000180",
        X"00000181",
        X"00000182",
        X"00000183",
        X"00000184",
        X"00000185",
        X"00000186",
        X"00000187",
        X"00000188",
        X"00000189",
        X"0000018a",
        X"0000018b",
        X"0000018c",
        X"0000018d",
        X"0000018e",
        X"0000018f",
        X"00000190",
        X"00000191",
        X"00000192",
        X"00000193",
        X"00000194",
        X"00000195",
        X"00000196",
        X"00000197",
        X"00000198",
        X"00000199",
        X"0000019a",
        X"0000019b",
        X"0000019c",
        X"0000019d",
        X"0000019e",
        X"0000019f",
        X"000001a0",
        X"000001a1",
        X"000001a2",
        X"000001a3",
        X"000001a4",
        X"000001a5",
        X"000001a6",
        X"000001a7",
        X"000001a8",
        X"000001a9",
        X"000001aa",
        X"000001ab",
        X"000001ac",
        X"000001ad",
        X"000001ae",
        X"000001af",
        X"000001b0",
        X"000001b1",
        X"000001b2",
        X"000001b3",
        X"000001b4",
        X"000001b5",
        X"000001b6",
        X"000001b7",
        X"000001b8",
        X"000001b9",
        X"000001ba",
        X"000001bb",
        X"000001bc",
        X"000001bd",
        X"000001be",
        X"000001bf",
        X"000001c0",
        X"000001c1",
        X"000001c2",
        X"000001c3",
        X"000001c4",
        X"000001c5",
        X"000001c6",
        X"000001c7",
        X"000001c8",
        X"000001c9",
        X"000001ca",
        X"000001cb",
        X"000001cc",
        X"000001cd",
        X"000001ce",
        X"000001cf",
        X"000001d0",
        X"000001d1",
        X"000001d2",
        X"000001d3",
        X"000001d4",
        X"000001d5",
        X"000001d6",
        X"000001d7",
        X"000001d8",
        X"000001d9",
        X"000001da",
        X"000001db",
        X"000001dc",
        X"000001dd",
        X"000001de",
        X"000001df",
        X"000001e0",
        X"000001e1",
        X"000001e2",
        X"000001e3",
        X"000001e4",
        X"000001e5",
        X"000001e6",
        X"000001e7",
        X"000001e8",
        X"000001e9",
        X"000001ea",
        X"000001eb",
        X"000001ec",
        X"000001ed",
        X"000001ee",
        X"000001ef",
        X"000001f0",
        X"000001f1",
        X"000001f2",
        X"000001f3",
        X"000001f4",
        X"000001f5",
        X"000001f6",
        X"000001f7",
        X"000001f8",
        X"000001f9",
        X"000001fa",
        X"000001fb",
        X"000001fc",
        X"000001fd",
        X"000001fe",
        X"000001ff",
        X"00000200",
        X"00000201",
        X"00000202",
        X"00000203",
        X"00000204",
        X"00000205",
        X"00000206",
        X"00000207",
        X"00000208",
        X"00000209",
        X"0000020a",
        X"0000020b",
        X"0000020c",
        X"0000020d",
        X"0000020e",
        X"0000020f",
        X"00000210",
        X"00000211",
        X"00000212",
        X"00000213",
        X"00000214",
        X"00000215",
        X"00000216",
        X"00000217",
        X"00000218",
        X"00000219",
        X"0000021a",
        X"0000021b",
        X"0000021c",
        X"0000021d",
        X"0000021e",
        X"0000021f",
        X"00000220",
        X"00000221",
        X"00000222",
        X"00000223",
        X"00000224",
        X"00000225",
        X"00000226",
        X"00000227",
        X"00000228",
        X"00000229",
        X"0000022a",
        X"0000022b",
        X"0000022c",
        X"0000022d",
        X"0000022e",
        X"0000022f",
        X"00000230",
        X"00000231",
        X"00000232",
        X"00000233",
        X"00000234",
        X"00000235",
        X"00000236",
        X"00000237",
        X"00000238",
        X"00000239",
        X"0000023a",
        X"0000023b",
        X"0000023c",
        X"0000023d",
        X"0000023e",
        X"0000023f",
        X"00000240",
        X"00000241",
        X"00000242",
        X"00000243",
        X"00000244",
        X"00000245",
        X"00000246",
        X"00000247",
        X"00000248",
        X"00000249",
        X"0000024a",
        X"0000024b",
        X"0000024c",
        X"0000024d",
        X"0000024e",
        X"0000024f",
        X"00000250",
        X"00000251",
        X"00000252",
        X"00000253",
        X"00000254",
        X"00000255",
        X"00000256",
        X"00000257",
        X"00000258",
        X"00000259",
        X"0000025a",
        X"0000025b",
        X"0000025c",
        X"0000025d",
        X"0000025e",
        X"0000025f",
        X"00000260",
        X"00000261",
        X"00000262",
        X"00000263",
        X"00000264",
        X"00000265",
        X"00000266",
        X"00000267",
        X"00000268",
        X"00000269",
        X"0000026a",
        X"0000026b",
        X"0000026c",
        X"0000026d",
        X"0000026e",
        X"0000026f",
        X"00000270",
        X"00000271",
        X"00000272",
        X"00000273",
        X"00000274",
        X"00000275",
        X"00000276",
        X"00000277",
        X"00000278",
        X"00000279",
        X"0000027a",
        X"0000027b",
        X"0000027c",
        X"0000027d",
        X"0000027e",
        X"0000027f",
        X"00000280",
        X"00000281",
        X"00000282",
        X"00000283",
        X"00000284",
        X"00000285",
        X"00000286",
        X"00000287",
        X"00000288",
        X"00000289",
        X"0000028a",
        X"0000028b",
        X"0000028c",
        X"0000028d",
        X"0000028e",
        X"0000028f",
        X"00000290",
        X"00000291",
        X"00000292",
        X"00000293",
        X"00000294",
        X"00000295",
        X"00000296",
        X"00000297",
        X"00000298",
        X"00000299",
        X"0000029a",
        X"0000029b",
        X"0000029c",
        X"0000029d",
        X"0000029e",
        X"0000029f",
        X"000002a0",
        X"000002a1",
        X"000002a2",
        X"000002a3",
        X"000002a4",
        X"000002a5",
        X"000002a6",
        X"000002a7",
        X"000002a8",
        X"000002a9",
        X"000002aa",
        X"000002ab",
        X"000002ac",
        X"000002ad",
        X"000002ae",
        X"000002af",
        X"000002b0",
        X"000002b1",
        X"000002b2",
        X"000002b3",
        X"000002b4",
        X"000002b5",
        X"000002b6",
        X"000002b7",
        X"000002b8",
        X"000002b9",
        X"000002ba",
        X"000002bb",
        X"000002bc",
        X"000002bd",
        X"000002be",
        X"000002bf",
        X"000002c0",
        X"000002c1",
        X"000002c2",
        X"000002c3",
        X"000002c4",
        X"000002c5",
        X"000002c6",
        X"000002c7",
        X"000002c8",
        X"000002c9",
        X"000002ca",
        X"000002cb",
        X"000002cc",
        X"000002cd",
        X"000002ce",
        X"000002cf",
        X"000002d0",
        X"000002d1",
        X"000002d2",
        X"000002d3",
        X"000002d4",
        X"000002d5",
        X"000002d6",
        X"000002d7",
        X"000002d8",
        X"000002d9",
        X"000002da",
        X"000002db",
        X"000002dc",
        X"000002dd",
        X"000002de",
        X"000002df",
        X"000002e0",
        X"000002e1",
        X"000002e2",
        X"000002e3",
        X"000002e4",
        X"000002e5",
        X"000002e6",
        X"000002e7",
        X"000002e8",
        X"000002e9",
        X"000002ea",
        X"000002eb",
        X"000002ec",
        X"000002ed",
        X"000002ee",
        X"000002ef",
        X"000002f0",
        X"000002f1",
        X"000002f2",
        X"000002f3",
        X"000002f4",
        X"000002f5",
        X"000002f6",
        X"000002f7",
        X"000002f8",
        X"000002f9",
        X"000002fa",
        X"000002fb",
        X"000002fc",
        X"000002fd",
        X"000002fe",
        X"000002ff",
        X"00000300",
        X"00000301",
        X"00000302",
        X"00000303",
        X"00000304",
        X"00000305",
        X"00000306",
        X"00000307",
        X"00000308",
        X"00000309",
        X"0000030a",
        X"0000030b",
        X"0000030c",
        X"0000030d",
        X"0000030e",
        X"0000030f",
        X"00000310",
        X"00000311",
        X"00000312",
        X"00000313",
        X"00000314",
        X"00000315",
        X"00000316",
        X"00000317",
        X"00000318",
        X"00000319",
        X"0000031a",
        X"0000031b",
        X"0000031c",
        X"0000031d",
        X"0000031e",
        X"0000031f",
        X"00000320",
        X"00000321",
        X"00000322",
        X"00000323",
        X"00000324",
        X"00000325",
        X"00000326",
        X"00000327",
        X"00000328",
        X"00000329",
        X"0000032a",
        X"0000032b",
        X"0000032c",
        X"0000032d",
        X"0000032e",
        X"0000032f",
        X"00000330",
        X"00000331",
        X"00000332",
        X"00000333",
        X"00000334",
        X"00000335",
        X"00000336",
        X"00000337",
        X"00000338",
        X"00000339",
        X"0000033a",
        X"0000033b",
        X"0000033c",
        X"0000033d",
        X"0000033e",
        X"0000033f",
        X"00000340",
        X"00000341",
        X"00000342",
        X"00000343",
        X"00000344",
        X"00000345",
        X"00000346",
        X"00000347",
        X"00000348",
        X"00000349",
        X"0000034a",
        X"0000034b",
        X"0000034c",
        X"0000034d",
        X"0000034e",
        X"0000034f",
        X"00000350",
        X"00000351",
        X"00000352",
        X"00000353",
        X"00000354",
        X"00000355",
        X"00000356",
        X"00000357",
        X"00000358",
        X"00000359",
        X"0000035a",
        X"0000035b",
        X"0000035c",
        X"0000035d",
        X"0000035e",
        X"0000035f",
        X"00000360",
        X"00000361",
        X"00000362",
        X"00000363",
        X"00000364",
        X"00000365",
        X"00000366",
        X"00000367",
        X"00000368",
        X"00000369",
        X"0000036a",
        X"0000036b",
        X"0000036c",
        X"0000036d",
        X"0000036e",
        X"0000036f",
        X"00000370",
        X"00000371",
        X"00000372",
        X"00000373",
        X"00000374",
        X"00000375",
        X"00000376",
        X"00000377",
        X"00000378",
        X"00000379",
        X"0000037a",
        X"0000037b",
        X"0000037c",
        X"0000037d",
        X"0000037e",
        X"0000037f",
        X"00000380",
        X"00000381",
        X"00000382",
        X"00000383",
        X"00000384",
        X"00000385",
        X"00000386",
        X"00000387",
        X"00000388",
        X"00000389",
        X"0000038a",
        X"0000038b",
        X"0000038c",
        X"0000038d",
        X"0000038e",
        X"0000038f",
        X"00000390",
        X"00000391",
        X"00000392",
        X"00000393",
        X"00000394",
        X"00000395",
        X"00000396",
        X"00000397",
        X"00000398",
        X"00000399",
        X"0000039a",
        X"0000039b",
        X"0000039c",
        X"0000039d",
        X"0000039e",
        X"0000039f",
        X"000003a0",
        X"000003a1",
        X"000003a2",
        X"000003a3",
        X"000003a4",
        X"000003a5",
        X"000003a6",
        X"000003a7",
        X"000003a8",
        X"000003a9",
        X"000003aa",
        X"000003ab",
        X"000003ac",
        X"000003ad",
        X"000003ae",
        X"000003af",
        X"000003b0",
        X"000003b1",
        X"000003b2",
        X"000003b3",
        X"000003b4",
        X"000003b5",
        X"000003b6",
        X"000003b7",
        X"000003b8",
        X"000003b9",
        X"000003ba",
        X"000003bb",
        X"000003bc",
        X"000003bd",
        X"000003be",
        X"000003bf",
        X"000003c0",
        X"000003c1",
        X"000003c2",
        X"000003c3",
        X"000003c4",
        X"000003c5",
        X"000003c6",
        X"000003c7",
        X"000003c8",
        X"000003c9",
        X"000003ca",
        X"000003cb",
        X"000003cc",
        X"000003cd",
        X"000003ce",
        X"000003cf",
        X"000003d0",
        X"000003d1",
        X"000003d2",
        X"000003d3",
        X"000003d4",
        X"000003d5",
        X"000003d6",
        X"000003d7",
        X"000003d8",
        X"000003d9",
        X"000003da",
        X"000003db",
        X"000003dc",
        X"000003dd",
        X"000003de",
        X"000003df",
        X"000003e0",
        X"000003e1",
        X"000003e2",
        X"000003e3",
        X"000003e4",
        X"000003e5",
        X"000003e6",
        X"000003e7",
        X"000003e8",
        X"000003e9",
        X"000003ea",
        X"000003eb",
        X"000003ec",
        X"000003ed",
        X"000003ee",
        X"000003ef",
        X"000003f0",
        X"000003f1",
        X"000003f2",
        X"000003f3",
        X"000003f4",
        X"000003f5",
        X"000003f6",
        X"000003f7",
        X"000003f8",
        X"000003f9",
        X"000003fa",
        X"000003fb",
        X"000003fc",
        X"000003fd",
        X"000003fe",
        X"000003ff"
    );

    attribute ram_style : string;
    attribute ram_style of table : signal is "block";

begin
    process (clk_i) begin
        if rising_edge(clk_i) then
            dat_o <= table(to_integer(addr_i));
        end if;
    end process;
end;
